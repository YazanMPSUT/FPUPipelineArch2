//`include "IPAdder.sv"
//`include "IMemory.sv"
//`include "Decode.sv"
//`include "RegisterFile.sv"
//`include "SetFlags.sv"
`include "Forward.sv"
`include "Buffer_IFID.sv"
`include "Buffer_IDEX.sv"
`include "Buffer_EXWB.sv"
`include "CommonClock.sv"
`include "MUX32.sv"
`include "EXE.sv"
`include "FetchStage.sv"
`include "DecodeStage.sv"
//`include "FPU.sv"
